`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:27:32 06/14/2012 
// Design Name: 
// Module Name:    reorder_queue
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description:
// Reorders downstream TLPs to output in increasing tag sequence. Input packets
// are stored in RAM and then read out when all previous sequence numbers have
// arrived and been read out. This module also provides the next available tag
// for the TX engine to use when sending memory request TLPs.
//
// Dependencies: 
// reorder_queue_input.v
// reorder_queue_output.v
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module reorder_queue #(
	parameter C_PCI_DATA_WIDTH = 9'd128,
	parameter C_NUM_CHNL = 4'd12,
	parameter C_MAX_READ_REQ_BYTES = 512,			// Max size of read requests (in bytes)
	parameter C_TAG_WIDTH = 5, 						// Number of outstanding requests 
	// Local parameters
	parameter C_PCI_DATA_WORD = C_PCI_DATA_WIDTH/32,
	parameter C_PCI_DATA_COUNT_WIDTH = clog2(C_PCI_DATA_WORD+1),
	parameter C_NUM_TAGS = 2**C_TAG_WIDTH,
	parameter C_DW_PER_TAG = C_MAX_READ_REQ_BYTES/4,
	parameter C_TAG_DW_COUNT_WIDTH = clog2s(C_DW_PER_TAG+1),
	parameter C_DATA_ADDR_STRIDE_WIDTH = clog2s(C_DW_PER_TAG/C_PCI_DATA_WORD), // div by C_PCI_DATA_WORD b/c there are C_PCI_DATA_WORD RAMs
	parameter C_DATA_ADDR_WIDTH = C_TAG_WIDTH + C_DATA_ADDR_STRIDE_WIDTH
)
(
	input CLK,														// Clock
	input RST,														// Synchronous reset
	input VALID,													// Valid input packet
	input [C_PCI_DATA_WIDTH-1:0] DATA,								// Input packet payload
	input [C_PCI_DATA_WORD-1:0] DATA_EN,							// Input packet payload data enable
	input [C_PCI_DATA_COUNT_WIDTH-1:0] DATA_EN_COUNT,				// Input packet payload data enable count
	input DONE,														// Input packet done
	input ERR,														// Input packet has error
	input [C_TAG_WIDTH-1:0] TAG,									// Input packet tag (external tag)

	input [5:0] INT_TAG,											// Internal tag to exchange with external
	input INT_TAG_VALID,											// High to signal tag exchange 
	output [C_TAG_WIDTH-1:0] EXT_TAG,								// External tag to provide in exchange for internal tag
	output EXT_TAG_VALID,											// High to signal external tag is valid

	output [C_PCI_DATA_WIDTH-1:0] ENG_DATA,							// Engine data 
	output [(C_NUM_CHNL*C_PCI_DATA_COUNT_WIDTH)-1:0] MAIN_DATA_EN,	// Main data enable
	output [C_NUM_CHNL-1:0] MAIN_DONE,								// Main data complete
	output [C_NUM_CHNL-1:0] MAIN_ERR,								// Main data completed with error
	output [(C_NUM_CHNL*C_PCI_DATA_COUNT_WIDTH)-1:0] SG_RX_DATA_EN,	// Scatter gather for RX data enable
	output [C_NUM_CHNL-1:0] SG_RX_DONE,								// Scatter gather for RX data complete
	output [C_NUM_CHNL-1:0] SG_RX_ERR,								// Scatter gather for RX data completed with error
	output [(C_NUM_CHNL*C_PCI_DATA_COUNT_WIDTH)-1:0] SG_TX_DATA_EN,	// Scatter gather for TX data enable
	output [C_NUM_CHNL-1:0] SG_TX_DONE,								// Scatter gather for TX data complete
	output [C_NUM_CHNL-1:0] SG_TX_ERR								// Scatter gather for TX data completed with error
);

`include "common_functions.v"

wire	[(C_DATA_ADDR_WIDTH*C_PCI_DATA_WORD)-1:0]	wWrDataAddr;
wire	[C_PCI_DATA_WIDTH-1:0]						wWrData;
wire	[C_PCI_DATA_WORD-1:0]						wWrDataEn;

wire	[C_TAG_WIDTH-1:0] 							wWrPktTag;
wire	[C_TAG_DW_COUNT_WIDTH-1:0] 					wWrPktWords;
wire							 					wWrPktWordsLTE1;
wire							 					wWrPktWordsLTE2;
wire							 					wWrPktValid;
wire							 					wWrPktDone;
wire							 					wWrPktErr;

wire	[C_DATA_ADDR_WIDTH-1:0]						wRdDataAddr;
wire	[C_PCI_DATA_WIDTH-1:0]						wRdData;

wire	[C_TAG_WIDTH-1:0] 							wRdPktTag;
wire	[(1+1+1+1+C_TAG_DW_COUNT_WIDTH)-1:0] 		wRdPktInfo;

wire	[5:0]										wRdTagMap;

reg		[C_TAG_WIDTH-1:0]							rPos=0;
reg													rValid=0;
wire	[C_NUM_TAGS-1:0]							wFinish;
reg		[C_NUM_TAGS-1:0]							rFinished=0;
reg		[C_NUM_TAGS-1:0]							rUse=0;
reg		[C_NUM_TAGS-1:0]							rUsing=0;
wire	[C_NUM_TAGS-1:0]							wClear;


assign EXT_TAG = rPos;
assign EXT_TAG_VALID = rValid;


// Move through tag/slot/bucket space.
always @ (posedge CLK) begin
	if (RST) begin
		rPos <= #1 0;
		rUse <= #1 0;
		rValid <= #1 0;
	end
	else begin
		if (INT_TAG_VALID & EXT_TAG_VALID) begin
			rPos <= #1 rPos + 1'd1;
			rUse <= #1 1<<rPos;
			rValid <= #1 !rUsing[rPos + 1'd1];
		end
		else begin
			rUse <= #1 0;
			rValid <= #1 !rUsing[rPos];
		end
	end
end


// Update tag/slot/bucket status.
always @ (posedge CLK) begin
	if (RST) begin
		rUsing <= #1 0;
		rFinished <= #1 0;
	end
	else begin
		rUsing <= #1 (rUsing | rUse) & ~wClear;
		rFinished <= #1 (rFinished | wFinish) & ~wClear;
	end
end


genvar r;
generate
	for (r = 0; r < C_PCI_DATA_WORD; r = r + 1) begin : rams
		// RAMs for packet reordering.
		(* RAM_STYLE="BLOCK" *)
		ram_1clk_1w_1r #(.C_RAM_WIDTH(32), .C_RAM_DEPTH(C_NUM_TAGS*C_DW_PER_TAG/C_PCI_DATA_WORD)) ram (
			.CLK(CLK),
			.ADDRA(wWrDataAddr[C_DATA_ADDR_WIDTH*r +:C_DATA_ADDR_WIDTH]),
			.WEA(wWrDataEn[r]),
			.DINA(wWrData[32*r +:32]),
			.ADDRB(wRdDataAddr),
			.DOUTB(wRdData[32*r +:32])
		);
	end
endgenerate


// RAM for bucket done, err, final DW count
(* RAM_STYLE="DISTRIBUTED" *)
ram_1clk_1w_1r #(.C_RAM_WIDTH(1 + 1 + 1 + 1 + C_TAG_DW_COUNT_WIDTH), .C_RAM_DEPTH(C_NUM_TAGS)) pktRam (
	.CLK(CLK),
	.ADDRA(wWrPktTag),
	.WEA((wWrPktDone | wWrPktErr) & wWrPktValid),
	.DINA({wWrPktDone, wWrPktErr, wWrPktWordsLTE2, wWrPktWordsLTE1, wWrPktWords}),
	.ADDRB(wRdPktTag),
	.DOUTB(wRdPktInfo)
);


// RAM for tag map
(* RAM_STYLE="DISTRIBUTED" *)
ram_1clk_1w_1r #(.C_RAM_WIDTH(6), .C_RAM_DEPTH(C_NUM_TAGS)) mapRam (
	.CLK(CLK),
	.ADDRA(rPos),
	.WEA(INT_TAG_VALID & EXT_TAG_VALID),
	.DINA(INT_TAG),
	.ADDRB(wRdPktTag),
	.DOUTB(wRdTagMap)
);


// Demux input data into the correct slot/bucket.
reorder_queue_input #(
	.C_PCI_DATA_WIDTH(C_PCI_DATA_WIDTH),
	.C_TAG_WIDTH(C_TAG_WIDTH),
	.C_TAG_DW_COUNT_WIDTH(C_TAG_DW_COUNT_WIDTH),
	.C_DATA_ADDR_STRIDE_WIDTH(C_DATA_ADDR_STRIDE_WIDTH),
	.C_DATA_ADDR_WIDTH(C_DATA_ADDR_WIDTH)
) data_input (
	.CLK(CLK),
	.RST(RST),
	.VALID(VALID),
	.DATA(DATA),
	.DATA_EN(DATA_EN),
	.DATA_EN_COUNT(DATA_EN_COUNT),
	.DONE(DONE),
	.ERR(ERR),
	.TAG(TAG),
	.TAG_FINISH(wFinish),
	.TAG_CLEAR(wClear),
	.STORED_DATA_ADDR(wWrDataAddr),
	.STORED_DATA(wWrData),
	.STORED_DATA_EN(wWrDataEn),
	.PKT_VALID(wWrPktValid),
	.PKT_TAG(wWrPktTag),
	.PKT_WORDS(wWrPktWords),
	.PKT_WORDS_LTE1(wWrPktWordsLTE1),
	.PKT_WORDS_LTE2(wWrPktWordsLTE2),
	.PKT_DONE(wWrPktDone),
	.PKT_ERR(wWrPktErr)
);


// Output packets in increasing tag order.
reorder_queue_output #(
	.C_PCI_DATA_WIDTH(C_PCI_DATA_WIDTH),
	.C_NUM_CHNL(C_NUM_CHNL),
	.C_TAG_WIDTH(C_TAG_WIDTH),
	.C_TAG_DW_COUNT_WIDTH(C_TAG_DW_COUNT_WIDTH),
	.C_DATA_ADDR_STRIDE_WIDTH(C_DATA_ADDR_STRIDE_WIDTH),
	.C_DATA_ADDR_WIDTH(C_DATA_ADDR_WIDTH)
) data_output (
	.CLK(CLK),
	.RST(RST),
	.DATA_ADDR(wRdDataAddr),
	.DATA(wRdData),
	.TAG_FINISHED(rFinished),
	.TAG_CLEAR(wClear),
	.TAG(wRdPktTag),
	.TAG_MAPPED(wRdTagMap),
	.PKT_WORDS(wRdPktInfo[0 +:C_TAG_DW_COUNT_WIDTH]),
	.PKT_WORDS_LTE1(wRdPktInfo[C_TAG_DW_COUNT_WIDTH]),
	.PKT_WORDS_LTE2(wRdPktInfo[C_TAG_DW_COUNT_WIDTH+1]),
	.PKT_ERR(wRdPktInfo[C_TAG_DW_COUNT_WIDTH+2]),
	.PKT_DONE(wRdPktInfo[C_TAG_DW_COUNT_WIDTH+3]),
	.ENG_DATA(ENG_DATA),
	.MAIN_DATA_EN(MAIN_DATA_EN),
	.MAIN_DONE(MAIN_DONE),
	.MAIN_ERR(MAIN_ERR),
	.SG_RX_DATA_EN(SG_RX_DATA_EN),
	.SG_RX_DONE(SG_RX_DONE),
	.SG_RX_ERR(SG_RX_ERR),
	.SG_TX_DATA_EN(SG_TX_DATA_EN),
	.SG_TX_DONE(SG_TX_DONE),
	.SG_TX_ERR(SG_TX_ERR)
);



/*
wire [35:0] wControl0;
chipscope_icon_1 cs_icon(
	.CONTROL0(wControl0)
);

chipscope_ila_t8_512_max a0(
	.CLK(CLK), 
	.CONTROL(wControl0), 
	.TRIG0({(MAIN_DATA_EN != 0 || MAIN_ERR != 0 || MAIN_DONE != 0 || SG_RX_DATA_EN != 0 || SG_RX_DONE != 0 || SG_RX_ERR != 0 || SG_TX_DATA_EN != 0 || SG_TX_DONE != 0 || SG_TX_ERR != 0),
		wWrDataEn != 0, wWrPktValid, wClear != 0, wFinish != 0, VALID, 2'd0}),
	.DATA({
			DATA[105:0], // 106
			SG_TX_ERR, // 2
			SG_TX_DONE, // 2
			SG_TX_DATA_EN, // 6
			SG_RX_ERR, // 2
			SG_RX_DONE, // 2
			SG_RX_DATA_EN, // 6
			MAIN_ERR, // 2
			MAIN_DONE, // 2
			MAIN_DATA_EN, // 6
			EXT_TAG_VALID, // 1
			INT_TAG_VALID, // 1
			TAG, // 5
			ERR, // 1
			DONE, // 1
			DATA_EN_COUNT, // 3
			DATA_EN, // 4
			VALID, // 1
			wWrDataAddr, // 40
			wWrData, // 128
			wWrDataEn, // 4
			wWrPktTag, // 5
			wWrPktWords, // 8
			wWrPktWordsLTE1, // 1
			wWrPktWordsLTE2, // 1
			wWrPktValid, // 1
			wWrPktDone, // 1
			wWrPktErr, // 1
			wRdDataAddr, // 10
			wRdPktTag, // 5
			wRdPktInfo, // 12
			wRdTagMap, // 6
			wFinish, // 32
			rFinished, // 32
			rUsing, // 32
			wClear, // 32
			rValid, // 1
			rPos, // 5
			2'd0}) // 2
);
*/

endmodule
